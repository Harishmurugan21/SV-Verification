Compiler version U-2023.03-SP2_Full64; Runtime version U-2023.03-SP2_Full64;  Dec 18 02:37 2025
generator class signal
$time=0| rst=0 | d=1 | q=0 |
generator class signal
$time=0| rst=1 | d=0 | q=0 |
generator class signal
$time=0| rst=0 | d=0 | q=0 |
generator class signal
$time=0| rst=1 | d=0 | q=0 |
generator class signal
$time=0| rst=0 | d=1 | q=0 |
generator class signal
$time=0| rst=0 | d=0 | q=0 |
generator class signal
$time=0| rst=1 | d=1 | q=0 |
generator class signal
$time=0| rst=1 | d=1 | q=0 |
generator class signal
$time=0| rst=0 | d=0 | q=0 |
generator class signal
$time=0| rst=1 | d=1 | q=0 |
generator class signal
$time=0| rst=0 | d=1 | q=0 |
generator class signal
$time=0| rst=0 | d=1 | q=0 |
generator class signal
$time=0| rst=1 | d=1 | q=0 |
generator class signal
$time=0| rst=0 | d=1 | q=0 |
generator class signal
$time=0| rst=1 | d=1 | q=0 |
------All sample testcases generated----------
monitor class signals
$time=6| rst=0 | d=0 | q=0 |
signals received on score board
$time=6| rst=0 | d=0 | q=0 |
-------pass--------
driver signal
$time=10| rst=0 | d=1 | q=0 |
monitor class signals
$time=16| rst=0 | d=1 | q=1 |
signals received on score board
$time=16| rst=0 | d=1 | q=1 |
-------pass--------
driver signal
$time=20| rst=1 | d=0 | q=0 |
monitor class signals
$time=26| rst=1 | d=1 | q=0 |
signals received on score board
$time=26| rst=1 | d=1 | q=0 |
-------pass--------
driver signal
$time=30| rst=0 | d=0 | q=0 |
monitor class signals
$time=36| rst=0 | d=0 | q=0 |
signals received on score board
$time=36| rst=0 | d=0 | q=0 |
-------pass--------
driver signal
$time=40| rst=1 | d=0 | q=0 |
monitor class signals
$time=46| rst=1 | d=0 | q=0 |
signals received on score board
$time=46| rst=1 | d=0 | q=0 |
-------pass--------
driver signal
$time=50| rst=0 | d=1 | q=0 |
monitor class signals
$time=56| rst=0 | d=1 | q=1 |
signals received on score board
$time=56| rst=0 | d=1 | q=1 |
-------pass--------
driver signal
$time=60| rst=0 | d=0 | q=0 |
monitor class signals
$time=66| rst=0 | d=0 | q=0 |
signals received on score board
$time=66| rst=0 | d=0 | q=0 |
-------pass--------
driver signal
$time=70| rst=1 | d=1 | q=0 |
monitor class signals
$time=76| rst=1 | d=0 | q=0 |
signals received on score board
$time=76| rst=1 | d=0 | q=0 |
-------pass--------
driver signal
$time=80| rst=1 | d=1 | q=0 |
monitor class signals
$time=86| rst=1 | d=0 | q=0 |
signals received on score board
$time=86| rst=1 | d=0 | q=0 |
-------pass--------
driver signal
$time=90| rst=0 | d=0 | q=0 |
monitor class signals
$time=96| rst=0 | d=0 | q=0 |
signals received on score board
$time=96| rst=0 | d=0 | q=0 |
-------pass--------
driver signal
$time=100| rst=1 | d=1 | q=0 |
monitor class signals
$time=106| rst=1 | d=0 | q=0 |
signals received on score board
$time=106| rst=1 | d=0 | q=0 |
-------pass--------
driver signal
$time=110| rst=0 | d=1 | q=0 |
monitor class signals
$time=116| rst=0 | d=1 | q=1 |
signals received on score board
$time=116| rst=0 | d=1 | q=1 |
-------pass--------
driver signal
$time=120| rst=0 | d=1 | q=0 |
monitor class signals
$time=126| rst=0 | d=1 | q=1 |
signals received on score board
$time=126| rst=0 | d=1 | q=1 |
-------pass--------
driver signal
$time=130| rst=1 | d=1 | q=0 |
monitor class signals
$time=136| rst=1 | d=1 | q=0 |
signals received on score board
$time=136| rst=1 | d=1 | q=0 |
-------pass--------
driver signal
$time=140| rst=0 | d=1 | q=0 |
monitor class signals
$time=146| rst=0 | d=1 | q=1 |
signals received on score board
$time=146| rst=0 | d=1 | q=1 |
-------pass--------
