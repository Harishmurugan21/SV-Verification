generator class signal
$time=0 | rst=0| w_en=0 | r_en=0 | data_in=00000000 |
generator class signal
$time=0 | rst=0| w_en=1 | r_en=0 | data_in=01101101 |
generator class signal
$time=0 | rst=0| w_en=1 | r_en=0 | data_in=11011101 |
generator class signal
$time=0 | rst=0| w_en=0 | r_en=0 | data_in=00000000 |
generator class signal
$time=0 | rst=0| w_en=1 | r_en=0 | data_in=00110010 |
generator class signal
$time=0 | rst=0| w_en=1 | r_en=0 | data_in=11011110 |
generator class signal
$time=0 | rst=0| w_en=1 | r_en=0 | data_in=00100110 |
generator class signal
$time=0 | rst=0| w_en=0 | r_en=0 | data_in=00000000 |
generator class signal
$time=0 | rst=0| w_en=1 | r_en=1 | data_in=00111000 |
generator class signal
$time=0 | rst=0| w_en=1 | r_en=0 | data_in=00110111 |
generator class signal
$time=0 | rst=0| w_en=1 | r_en=0 | data_in=00000111 |
generator class signal
$time=0 | rst=0| w_en=1 | r_en=1 | data_in=00011001 |
generator class signal
$time=0 | rst=0| w_en=1 | r_en=0 | data_in=10010100 |
generator class signal
$time=0 | rst=0| w_en=1 | r_en=0 | data_in=11010100 |
generator class signal
$time=0 | rst=0| w_en=1 | r_en=0 | data_in=10000010 |
generator class signal
$time=0 | rst=0| w_en=1 | r_en=0 | data_in=00110110 |
generator class signal
$time=0 | rst=0| w_en=1 | r_en=0 | data_in=11001110 |
generator class signal
$time=0 | rst=0| w_en=1 | r_en=1 | data_in=11010100 |
generator class signal
$time=0 | rst=0| w_en=1 | r_en=0 | data_in=11110111 |
generator class signal
$time=0 | rst=0| w_en=0 | r_en=0 | data_in=00000000 |
generator class signal
$time=0 | rst=0| w_en=1 | r_en=1 | data_in=01111000 |
generator class signal
$time=0 | rst=0| w_en=1 | r_en=0 | data_in=11110011 |
generator class signal
$time=0 | rst=0| w_en=1 | r_en=0 | data_in=10110001 |
generator class signal
$time=0 | rst=0| w_en=1 | r_en=0 | data_in=11110010 |
generator class signal
$time=0 | rst=0| w_en=1 | r_en=0 | data_in=00011000 |
generator class signal
$time=0 | rst=0| w_en=1 | r_en=0 | data_in=00101110 |
generator class signal
$time=0 | rst=0| w_en=1 | r_en=0 | data_in=01011111 |
generator class signal
$time=0 | rst=0| w_en=1 | r_en=1 | data_in=11110110 |
generator class signal
$time=0 | rst=0| w_en=1 | r_en=0 | data_in=00010011 |
generator class signal
$time=0 | rst=0| w_en=1 | r_en=1 | data_in=01010000 |
generator class signal
$time=0 | rst=0| w_en=1 | r_en=0 | data_in=10000100 |
generator class signal
$time=0 | rst=0| w_en=1 | r_en=0 | data_in=01001111 |
generator class signal
$time=0 | rst=0| w_en=1 | r_en=0 | data_in=01010110 |
generator class signal
$time=0 | rst=0| w_en=1 | r_en=0 | data_in=11000100 |
generator class signal
$time=0 | rst=0| w_en=1 | r_en=0 | data_in=10100010 |
generator class signal
$time=0 | rst=0| w_en=1 | r_en=0 | data_in=01100010 |
generator class signal
$time=0 | rst=0| w_en=1 | r_en=0 | data_in=00011100 |
generator class signal
$time=0 | rst=0| w_en=1 | r_en=0 | data_in=11101010 |
generator class signal
$time=0 | rst=0| w_en=1 | r_en=0 | data_in=00101101 |
generator class signal
$time=0 | rst=0| w_en=0 | r_en=0 | data_in=00000000 |
monitor class signals
$time=6 | rst=1| w_en=0 | r_en=0 | data_in=00000000 |data_out=00000000 | empty=1|full=0 | 
signals received on score board
$time=6 | rst=1| w_en=0 | r_en=0 | data_in=00000000 |data_out=00000000 | empty=1|full=0 | 
-------------------------------------------------
monitor class signals
$time=16 | rst=1| w_en=0 | r_en=0 | data_in=00000000 |data_out=00000000 | empty=1|full=0 | 
signals received on score board
$time=16 | rst=1| w_en=0 | r_en=0 | data_in=00000000 |data_out=00000000 | empty=1|full=0 | 
-------------------------------------------------
driver signal
$time=20 | rst=0| w_en=0 | r_en=0 | data_in=00000000 |
monitor class signals
$time=26 | rst=0| w_en=0 | r_en=0 | data_in=00000000 |data_out=00000000 | empty=1|full=0 | 
signals received on score board
$time=26 | rst=0| w_en=0 | r_en=0 | data_in=00000000 |data_out=00000000 | empty=1|full=0 | 
-------------------------------------------------
driver signal
$time=30 | rst=0| w_en=1 | r_en=0 | data_in=01101101 |
monitor class signals
$time=36 | rst=0| w_en=1 | r_en=0 | data_in=01101101 |data_out=00000000 | empty=0|full=0 | 
signals received on score board
$time=36 | rst=0| w_en=1 | r_en=0 | data_in=01101101 |data_out=00000000 | empty=0|full=0 | 
-------------------------------------------------
driver signal
$time=40 | rst=0| w_en=1 | r_en=0 | data_in=11011101 |
monitor class signals
$time=46 | rst=0| w_en=1 | r_en=0 | data_in=11011101 |data_out=00000000 | empty=0|full=0 | 
signals received on score board
$time=46 | rst=0| w_en=1 | r_en=0 | data_in=11011101 |data_out=00000000 | empty=0|full=0 | 
-------------------------------------------------
driver signal
$time=50 | rst=0| w_en=0 | r_en=0 | data_in=00000000 |
monitor class signals
$time=56 | rst=0| w_en=0 | r_en=0 | data_in=00000000 |data_out=00000000 | empty=0|full=0 | 
signals received on score board
$time=56 | rst=0| w_en=0 | r_en=0 | data_in=00000000 |data_out=00000000 | empty=0|full=0 | 
-------------------------------------------------
driver signal
$time=60 | rst=0| w_en=1 | r_en=0 | data_in=00110010 |
monitor class signals
$time=66 | rst=0| w_en=1 | r_en=0 | data_in=00110010 |data_out=00000000 | empty=0|full=0 | 
signals received on score board
$time=66 | rst=0| w_en=1 | r_en=0 | data_in=00110010 |data_out=00000000 | empty=0|full=0 | 
-------------------------------------------------
driver signal
$time=70 | rst=0| w_en=1 | r_en=0 | data_in=11011110 |
monitor class signals
$time=76 | rst=0| w_en=1 | r_en=0 | data_in=11011110 |data_out=00000000 | empty=0|full=0 | 
signals received on score board
$time=76 | rst=0| w_en=1 | r_en=0 | data_in=11011110 |data_out=00000000 | empty=0|full=0 | 
-------------------------------------------------
driver signal
$time=80 | rst=0| w_en=1 | r_en=0 | data_in=00100110 |
monitor class signals
$time=86 | rst=0| w_en=1 | r_en=0 | data_in=00100110 |data_out=00000000 | empty=0|full=0 | 
signals received on score board
$time=86 | rst=0| w_en=1 | r_en=0 | data_in=00100110 |data_out=00000000 | empty=0|full=0 | 
-------------------------------------------------
driver signal
$time=90 | rst=0| w_en=0 | r_en=0 | data_in=00000000 |
monitor class signals
$time=96 | rst=0| w_en=0 | r_en=0 | data_in=00000000 |data_out=00000000 | empty=0|full=0 | 
signals received on score board
$time=96 | rst=0| w_en=0 | r_en=0 | data_in=00000000 |data_out=00000000 | empty=0|full=0 | 
-------------------------------------------------
driver signal
$time=100 | rst=0| w_en=1 | r_en=1 | data_in=00111000 |
monitor class signals
$time=106 | rst=0| w_en=1 | r_en=1 | data_in=00111000 |data_out=01101101 | empty=0|full=0 | 
signals received on score board
$time=106 | rst=0| w_en=1 | r_en=1 | data_in=00111000 |data_out=01101101 | empty=0|full=0 | 
<---------pass--------->
-------------------------------------------------
driver signal
$time=110 | rst=0| w_en=1 | r_en=0 | data_in=00110111 |
monitor class signals
$time=116 | rst=0| w_en=1 | r_en=0 | data_in=00110111 |data_out=01101101 | empty=0|full=0 | 
signals received on score board
$time=116 | rst=0| w_en=1 | r_en=0 | data_in=00110111 |data_out=01101101 | empty=0|full=0 | 
-------------------------------------------------
driver signal
$time=120 | rst=0| w_en=1 | r_en=0 | data_in=00000111 |
monitor class signals
$time=126 | rst=0| w_en=1 | r_en=0 | data_in=00000111 |data_out=01101101 | empty=0|full=1 | 
signals received on score board
$time=126 | rst=0| w_en=1 | r_en=0 | data_in=00000111 |data_out=01101101 | empty=0|full=1 | 
-------------------------------------------------
driver signal
$time=130 | rst=0| w_en=1 | r_en=1 | data_in=00011001 |
monitor class signals
$time=136 | rst=0| w_en=1 | r_en=1 | data_in=00011001 |data_out=11011101 | empty=0|full=0 | 
signals received on score board
$time=136 | rst=0| w_en=1 | r_en=1 | data_in=00011001 |data_out=11011101 | empty=0|full=0 | 
<---------pass--------->
-------------------------------------------------
driver signal
$time=140 | rst=0| w_en=1 | r_en=0 | data_in=10010100 |
monitor class signals
$time=146 | rst=0| w_en=1 | r_en=0 | data_in=10010100 |data_out=11011101 | empty=0|full=1 | 
signals received on score board
$time=146 | rst=0| w_en=1 | r_en=0 | data_in=10010100 |data_out=11011101 | empty=0|full=1 | 
-------------------------------------------------
driver signal
$time=150 | rst=0| w_en=1 | r_en=0 | data_in=11010100 |
monitor class signals
$time=156 | rst=0| w_en=1 | r_en=0 | data_in=11010100 |data_out=11011101 | empty=0|full=1 | 
signals received on score board
$time=156 | rst=0| w_en=1 | r_en=0 | data_in=11010100 |data_out=11011101 | empty=0|full=1 | 
-------------------------------------------------
driver signal
$time=160 | rst=0| w_en=1 | r_en=0 | data_in=10000010 |
monitor class signals
$time=166 | rst=0| w_en=1 | r_en=0 | data_in=10000010 |data_out=11011101 | empty=0|full=1 | 
signals received on score board
$time=166 | rst=0| w_en=1 | r_en=0 | data_in=10000010 |data_out=11011101 | empty=0|full=1 | 
-------------------------------------------------
driver signal
$time=170 | rst=0| w_en=1 | r_en=0 | data_in=00110110 |
monitor class signals
$time=176 | rst=0| w_en=1 | r_en=0 | data_in=00110110 |data_out=11011101 | empty=0|full=1 | 
signals received on score board
$time=176 | rst=0| w_en=1 | r_en=0 | data_in=00110110 |data_out=11011101 | empty=0|full=1 | 
-------------------------------------------------
driver signal
$time=180 | rst=0| w_en=1 | r_en=0 | data_in=11001110 |
monitor class signals
$time=186 | rst=0| w_en=1 | r_en=0 | data_in=11001110 |data_out=11011101 | empty=0|full=1 | 
signals received on score board
$time=186 | rst=0| w_en=1 | r_en=0 | data_in=11001110 |data_out=11011101 | empty=0|full=1 | 
-------------------------------------------------
driver signal
$time=190 | rst=0| w_en=1 | r_en=1 | data_in=11010100 |
monitor class signals
$time=196 | rst=0| w_en=1 | r_en=1 | data_in=11010100 |data_out=00110010 | empty=0|full=0 | 
signals received on score board
$time=196 | rst=0| w_en=1 | r_en=1 | data_in=11010100 |data_out=00110010 | empty=0|full=0 | 
<---------pass--------->
-------------------------------------------------
driver signal
$time=200 | rst=0| w_en=1 | r_en=0 | data_in=11110111 |
monitor class signals
$time=206 | rst=0| w_en=1 | r_en=0 | data_in=11110111 |data_out=00110010 | empty=0|full=1 | 
signals received on score board
$time=206 | rst=0| w_en=1 | r_en=0 | data_in=11110111 |data_out=00110010 | empty=0|full=1 | 
-------------------------------------------------
driver signal
$time=210 | rst=0| w_en=0 | r_en=0 | data_in=00000000 |
monitor class signals
$time=216 | rst=0| w_en=0 | r_en=0 | data_in=00000000 |data_out=00110010 | empty=0|full=1 | 
signals received on score board
$time=216 | rst=0| w_en=0 | r_en=0 | data_in=00000000 |data_out=00110010 | empty=0|full=1 | 
-------------------------------------------------
driver signal
$time=220 | rst=0| w_en=1 | r_en=1 | data_in=01111000 |
monitor class signals
$time=226 | rst=0| w_en=1 | r_en=1 | data_in=01111000 |data_out=11011110 | empty=0|full=0 | 
signals received on score board
$time=226 | rst=0| w_en=1 | r_en=1 | data_in=01111000 |data_out=11011110 | empty=0|full=0 | 
<---------pass--------->
-------------------------------------------------
driver signal
$time=230 | rst=0| w_en=1 | r_en=0 | data_in=11110011 |
monitor class signals
$time=236 | rst=0| w_en=1 | r_en=0 | data_in=11110011 |data_out=11011110 | empty=0|full=1 | 
signals received on score board
$time=236 | rst=0| w_en=1 | r_en=0 | data_in=11110011 |data_out=11011110 | empty=0|full=1 | 
-------------------------------------------------
driver signal
$time=240 | rst=0| w_en=1 | r_en=0 | data_in=10110001 |
monitor class signals
$time=246 | rst=0| w_en=1 | r_en=0 | data_in=10110001 |data_out=11011110 | empty=0|full=1 | 
signals received on score board
$time=246 | rst=0| w_en=1 | r_en=0 | data_in=10110001 |data_out=11011110 | empty=0|full=1 | 
-------------------------------------------------
driver signal
$time=250 | rst=0| w_en=1 | r_en=0 | data_in=11110010 |
monitor class signals
$time=256 | rst=0| w_en=1 | r_en=0 | data_in=11110010 |data_out=11011110 | empty=0|full=1 | 
signals received on score board
$time=256 | rst=0| w_en=1 | r_en=0 | data_in=11110010 |data_out=11011110 | empty=0|full=1 | 
-------------------------------------------------
driver signal
$time=260 | rst=0| w_en=1 | r_en=0 | data_in=00011000 |
monitor class signals
$time=266 | rst=0| w_en=1 | r_en=0 | data_in=00011000 |data_out=11011110 | empty=0|full=1 | 
signals received on score board
$time=266 | rst=0| w_en=1 | r_en=0 | data_in=00011000 |data_out=11011110 | empty=0|full=1 | 
-------------------------------------------------
driver signal
$time=270 | rst=0| w_en=1 | r_en=0 | data_in=00101110 |
monitor class signals
$time=276 | rst=0| w_en=1 | r_en=0 | data_in=00101110 |data_out=11011110 | empty=0|full=1 | 
signals received on score board
$time=276 | rst=0| w_en=1 | r_en=0 | data_in=00101110 |data_out=11011110 | empty=0|full=1 | 
-------------------------------------------------
driver signal
$time=280 | rst=0| w_en=1 | r_en=0 | data_in=01011111 |
monitor class signals
$time=286 | rst=0| w_en=1 | r_en=0 | data_in=01011111 |data_out=11011110 | empty=0|full=1 | 
signals received on score board
$time=286 | rst=0| w_en=1 | r_en=0 | data_in=01011111 |data_out=11011110 | empty=0|full=1 | 
-------------------------------------------------
driver signal
$time=290 | rst=0| w_en=1 | r_en=1 | data_in=11110110 |
monitor class signals
$time=296 | rst=0| w_en=1 | r_en=1 | data_in=11110110 |data_out=00100110 | empty=0|full=0 | 
signals received on score board
$time=296 | rst=0| w_en=1 | r_en=1 | data_in=11110110 |data_out=00100110 | empty=0|full=0 | 
<---------pass--------->
-------------------------------------------------
driver signal
$time=300 | rst=0| w_en=1 | r_en=0 | data_in=00010011 |
monitor class signals
$time=306 | rst=0| w_en=1 | r_en=0 | data_in=00010011 |data_out=00100110 | empty=0|full=1 | 
signals received on score board
$time=306 | rst=0| w_en=1 | r_en=0 | data_in=00010011 |data_out=00100110 | empty=0|full=1 | 
-------------------------------------------------
driver signal
$time=310 | rst=0| w_en=1 | r_en=1 | data_in=01010000 |
monitor class signals
$time=316 | rst=0| w_en=1 | r_en=1 | data_in=01010000 |data_out=00111000 | empty=0|full=0 | 
signals received on score board
$time=316 | rst=0| w_en=1 | r_en=1 | data_in=01010000 |data_out=00111000 | empty=0|full=0 | 
<---------pass--------->
-------------------------------------------------
driver signal
$time=320 | rst=0| w_en=1 | r_en=0 | data_in=10000100 |
monitor class signals
$time=326 | rst=0| w_en=1 | r_en=0 | data_in=10000100 |data_out=00111000 | empty=0|full=1 | 
signals received on score board
$time=326 | rst=0| w_en=1 | r_en=0 | data_in=10000100 |data_out=00111000 | empty=0|full=1 | 
-------------------------------------------------
driver signal
$time=330 | rst=0| w_en=1 | r_en=0 | data_in=01001111 |
monitor class signals
$time=336 | rst=0| w_en=1 | r_en=0 | data_in=01001111 |data_out=00111000 | empty=0|full=1 | 
signals received on score board
$time=336 | rst=0| w_en=1 | r_en=0 | data_in=01001111 |data_out=00111000 | empty=0|full=1 | 
-------------------------------------------------
driver signal
$time=340 | rst=0| w_en=1 | r_en=0 | data_in=01010110 |
monitor class signals
$time=346 | rst=0| w_en=1 | r_en=0 | data_in=01010110 |data_out=00111000 | empty=0|full=1 | 
signals received on score board
$time=346 | rst=0| w_en=1 | r_en=0 | data_in=01010110 |data_out=00111000 | empty=0|full=1 | 
-------------------------------------------------
driver signal
$time=350 | rst=0| w_en=1 | r_en=0 | data_in=11000100 |
monitor class signals
$time=356 | rst=0| w_en=1 | r_en=0 | data_in=11000100 |data_out=00111000 | empty=0|full=1 | 
signals received on score board
$time=356 | rst=0| w_en=1 | r_en=0 | data_in=11000100 |data_out=00111000 | empty=0|full=1 | 
-------------------------------------------------
driver signal
$time=360 | rst=0| w_en=1 | r_en=0 | data_in=10100010 |
monitor class signals
$time=366 | rst=0| w_en=1 | r_en=0 | data_in=10100010 |data_out=00111000 | empty=0|full=1 | 
signals received on score board
$time=366 | rst=0| w_en=1 | r_en=0 | data_in=10100010 |data_out=00111000 | empty=0|full=1 | 
-------------------------------------------------
driver signal
$time=370 | rst=0| w_en=1 | r_en=0 | data_in=01100010 |
monitor class signals
$time=376 | rst=0| w_en=1 | r_en=0 | data_in=01100010 |data_out=00111000 | empty=0|full=1 | 
signals received on score board
$time=376 | rst=0| w_en=1 | r_en=0 | data_in=01100010 |data_out=00111000 | empty=0|full=1 | 
-------------------------------------------------
driver signal
$time=380 | rst=0| w_en=1 | r_en=0 | data_in=00011100 |
monitor class signals
$time=386 | rst=0| w_en=1 | r_en=0 | data_in=00011100 |data_out=00111000 | empty=0|full=1 | 
signals received on score board
$time=386 | rst=0| w_en=1 | r_en=0 | data_in=00011100 |data_out=00111000 | empty=0|full=1 | 
-------------------------------------------------
driver signal
$time=390 | rst=0| w_en=1 | r_en=0 | data_in=11101010 |
monitor class signals
$time=396 | rst=0| w_en=1 | r_en=0 | data_in=11101010 |data_out=00111000 | empty=0|full=1 | 
signals received on score board
$time=396 | rst=0| w_en=1 | r_en=0 | data_in=11101010 |data_out=00111000 | empty=0|full=1 | 
-------------------------------------------------
driver signal
$time=400 | rst=0| w_en=1 | r_en=0 | data_in=00101101 |
driver signal
$time=410 | rst=0| w_en=0 | r_en=0 | data_in=00000000 |
$finish called from file "testbench.sv", line 40.
$finish at simulation time                  600
