Compiler version U-2023.03-SP2_Full64; Runtime version U-2023.03-SP2_Full64;  Dec 22 13:34 2025
generatd class signal
time=0|rst=0| en=1| q=xxxxxx|
generatd class signal
time=0|rst=0| en=1| q=xxxxxx|
generatd class signal
time=0|rst=0| en=1| q=xxxxxx|
generatd class signal
time=0|rst=0| en=1| q=xxxxxx|
generatd class signal
time=0|rst=0| en=1| q=xxxxxx|
generatd class signal
time=0|rst=0| en=1| q=xxxxxx|
generatd class signal
time=0|rst=0| en=1| q=xxxxxx|
generatd class signal
time=0|rst=0| en=1| q=xxxxxx|
generatd class signal
time=0|rst=0| en=1| q=xxxxxx|
generatd class signal
time=0|rst=0| en=1| q=xxxxxx|
-------------------------------------------
monitor class signals
time=6|rst=1|en=0| q=0|
signals received on score board
time=6|rst=1|en=0| q=0|
----------pass---------
-------------------------------------------------
monitor class signals
time=16|rst=1|en=0| q=0|
signals received on score board
time=16|rst=1|en=0| q=0|
----------pass---------
-------------------------------------------------
driver class signal
time=20|rst=0| en=1| q=xxxxxx|
monitor class signals
time=26|rst=0| en=1| q=1|
signals received on score board
time=26|rst=0| en=1| q=1|
----------pass---------
-------------------------------------------------
driver class signal
time=30|rst=0| en=1| q=xxxxxx|
monitor class signals
time=36|rst=0| en=1| q=10|
signals received on score board
time=36|rst=0| en=1| q=10|
----------pass---------
-------------------------------------------------
driver class signal
time=40|rst=0| en=1| q=xxxxxx|
monitor class signals
time=46|rst=0| en=1| q=11|
signals received on score board
time=46|rst=0| en=1| q=11|
----------pass---------
-------------------------------------------------
driver class signal
time=50|rst=0| en=1| q=xxxxxx|
monitor class signals
time=56|rst=0| en=1| q=100|
signals received on score board
time=56|rst=0| en=1| q=100|
----------pass---------
-------------------------------------------------
driver class signal
time=60|rst=0| en=1| q=xxxxxx|
monitor class signals
time=66|rst=0| en=1| q=101|
signals received on score board
time=66|rst=0| en=1| q=101|
----------pass---------
-------------------------------------------------
driver class signal
time=70|rst=0| en=1| q=xxxxxx|
monitor class signals
time=76|rst=0| en=1| q=110|
signals received on score board
time=76|rst=0| en=1| q=110|
----------pass---------
-------------------------------------------------
driver class signal
time=80|rst=0| en=1| q=xxxxxx|
monitor class signals
time=86|rst=0| en=1| q=111|
signals received on score board
time=86|rst=0| en=1| q=111|
----------pass---------
-------------------------------------------------
driver class signal
time=90|rst=0| en=1| q=xxxxxx|
monitor class signals
time=96|rst=0| en=1| q=1000|
signals received on score board
time=96|rst=0| en=1| q=1000|
----------pass---------
-------------------------------------------------
driver class signal
time=100|rst=0| en=1| q=xxxxxx|
monitor class signals
time=106|rst=0| en=1| q=1001|
signals received on score board
time=106|rst=0| en=1| q=1001|
----------pass---------
-------------------------------------------------
driver class signal
time=110|rst=0| en=1| q=xxxxxx|
monitor class signals
time=116|rst=0| en=1| q=1010|
signals received on score board
time=116|rst=0| en=1| q=1010|
----------pass---------
-------------------------------------------------
$finish called from file "testbench.sv", 
